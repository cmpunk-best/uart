---
--UART main file for entity and architecture
---
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity main is
  port (
	--TODO
  ) ;
end entity ; -- main

architecture struct of main is

	signal 

begin
--TODO
end architecture ; -- struct